#Creates a directory for your project called "test" in your user directory
mkdir ~/git/test 
# Changes the current working directory to your newly created directory
cd ~/git/test

# Sets up the necessary Git files
git init
# Initialized empty Git repository in /Users/you/Hello-World/.git/

#Creates a file called "README.sv" in gitHub
##Creates a file called "README.loc" in gitHub
